interface crc7_if;
  logic sig_clk;
  logic sig_rst;
  logic sig_data;
  
  logic [6:0] sig_crc;
endinterface: crc7_if
